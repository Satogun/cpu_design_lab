module IF(


);


endmodule